`timescale 1ns/1ps

/* 

    * Assignment - 6
    * Problem - 3
    * Semester - 5 (Autumn)
    * Group - 56
    * Group members - Utsav Mehta (20CS10069) and Vibhu (20CS10072)

*/

module diff(a, b, out_diff);

    input [31:0] a, b;
    output reg [5:0] out_diff;

    wire [31:0] result, n, temp1, temp2;

    wire temp;
    assign n = a ^ b;
    
    adder_32_bit n_minus_one(.a(n), .b(32'b11111111111111111111111111111111), .c_in(1'b0), .sum(temp1), .c_out(temp));
    assign temp2 = temp1 ^ n;
    assign result = temp2 & n;

    // assign out_diff[5] = (a==b);

    always @(a, b) begin
        case (result)
            32'b00000000000000000000000000000000: out_diff[4:0] = 5'b00000;
            32'b00000000000000000000000000000001: out_diff[4:0] = 5'b00001;
            32'b00000000000000000000000000000010: out_diff[4:0] = 5'b00010;
            32'b00000000000000000000000000000100: out_diff[4:0] = 5'b00011;
            32'b00000000000000000000000000001000: out_diff[4:0] = 5'b00100;
            32'b00000000000000000000000000010000: out_diff[4:0] = 5'b00101;
            32'b00000000000000000000000000100000: out_diff[4:0] = 5'b00110;
            32'b00000000000000000000000001000000: out_diff[4:0] = 5'b00111;
            32'b00000000000000000000000010000000: out_diff[4:0] = 5'b01000;
            32'b00000000000000000000000100000000: out_diff[4:0] = 5'b01001;
            32'b00000000000000000000001000000000: out_diff[4:0] = 5'b01010;
            32'b00000000000000000000010000000000: out_diff[4:0] = 5'b01011;
            32'b00000000000000000000100000000000: out_diff[4:0] = 5'b01100;
            32'b00000000000000000001000000000000: out_diff[4:0] = 5'b01101;
            32'b00000000000000000010000000000000: out_diff[4:0] = 5'b01110;
            32'b00000000000000000100000000000000: out_diff[4:0] = 5'b01111;
            32'b00000000000000001000000000000000: out_diff[4:0] = 5'b10000;
            32'b00000000000000010000000000000000: out_diff[4:0] = 5'b10001;
            32'b00000000000000100000000000000000: out_diff[4:0] = 5'b10010;
            32'b00000000000001000000000000000000: out_diff[4:0] = 5'b10011;
            32'b00000000000010000000000000000000: out_diff[4:0] = 5'b10100;
            32'b00000000000100000000000000000000: out_diff[4:0] = 5'b10101;
            32'b00000000001000000000000000000000: out_diff[4:0] = 5'b10110;
            32'b00000000010000000000000000000000: out_diff[4:0] = 5'b10111;
            32'b00000000100000000000000000000000: out_diff[4:0] = 5'b11000;
            32'b00000001000000000000000000000000: out_diff[4:0] = 5'b11001;
            32'b00000010000000000000000000000000: out_diff[4:0] = 5'b11010;
            32'b00000100000000000000000000000000: out_diff[4:0] = 5'b11011;
            32'b00001000000000000000000000000000: out_diff[4:0] = 5'b11100;
            32'b00010000000000000000000000000000: out_diff[4:0] = 5'b11101;
            32'b00100000000000000000000000000000: out_diff[4:0] = 5'b11110;
            32'b01000000000000000000000000000000: out_diff[4:0] = 5'b11111;
            default: out_diff[4:0] = 5'b11111;
        endcase
    end
    
endmodule